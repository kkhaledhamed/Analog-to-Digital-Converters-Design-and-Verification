** sch_path: /home/tare/sar_adc/inv.sch
**.subckt inv Y A
*.ipin A
*.opin Y
**** begin user architecture code


*inverter model
a1 A Yi my_inv
.model my_inv d_inverter(rise_delay = 1e-9 fall_delay = 1e-9
+                        input_load = 1e-12)
*force netlisting of digital outputs
v1 Yi Y 0



.include /home/tare/pdk/gf180mcuC/libs.tech/ngspice/design.ngspice
.lib /home/tare/pdk/gf180mcuC/libs.tech/ngspice/sm141064.ngspice typical

**** end user architecture code
**.ends
.end
