** sch_path: /home/tare/Documents/sar_adc/inv_tb.sch
**.subckt inv_tb
V1 A GND pulse(0 VDD 0 TRF TRF {TCLK/2} {TCLK})
x1 Y A inv
**** begin user architecture code


*parameters
.param VDD=2 VCC=VDD
.param TRF=1n TCLK=100n
.param TSTOP={4*TCLK} TDROP=0

*analysis setup and control statements
.tran 1n {TSTOP} {TDROP}

*save all voltages and currents
.save all



.include /home/tare/pdk/gf180mcuC/libs.tech/ngspice/design.ngspice
.lib /home/tare/pdk/gf180mcuC/libs.tech/ngspice/sm141064.ngspice typical

**** end user architecture code
**.ends

* expanding   symbol:  /home/tare/Documents/sar_adc/inv.sym # of pins=2
** sym_path: /home/tare/Documents/sar_adc/inv.sym
** sch_path: /home/tare/Documents/sar_adc/inv.sch
.subckt inv Y A
*.ipin A
*.opin Y
**** begin user architecture code


*inverter model
a1 A Yi my_inv
.model my_inv d_inverter(rise_delay = 1e-9 fall_delay = 1e-9
+                        input_load = 1e-12)

*force netlisting of digital outputs
v1 Yi Y 0


**** end user architecture code
.ends

.GLOBAL GND
.end
